module sevenseg(output logic [6:0] hex_out, 
                input logic [3:0] data_in);

always_comb
  unique casez (data_in)
    4'b0000 : hex_out = 7'b1000000;
    4'b0001 : hex_out = 7'b1111001;
    4'b0010 : hex_out = 7'b0100100;
    4'b0011 : hex_out = 7'b0110000;
    4'b0100 : hex_out = 7'b0011001;
    4'b0101 : hex_out = 7'b0010010;
    4'b0110 : hex_out = 7'b0000010;
    4'b0111 : hex_out = 7'b1111000;
    4'b1000 : hex_out = 7'b0000000;
    4'b1001 : hex_out = 7'b0010000;
    4'b1010 : hex_out = 7'b0001000;
    4'b1011 : hex_out = 7'b0000011;
    4'b1100 : hex_out = 7'b1000110;
    4'b1101 : hex_out = 7'b0100001;
    4'b1110 : hex_out = 7'b0000110;
    4'b1111 : hex_out = 7'b0001110;
    default : hex_out = 7'b1111111;
  endcase
endmodule